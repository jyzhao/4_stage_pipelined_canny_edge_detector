library verilog;
use verilog.vl_types.all;
entity tb_gradient_magnitude_wrapper is
end tb_gradient_magnitude_wrapper;
