library verilog;
use verilog.vl_types.all;
entity tb_pts_sr is
end tb_pts_sr;
