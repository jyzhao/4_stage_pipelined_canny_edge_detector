library verilog;
use verilog.vl_types.all;
entity tb_gradient is
end tb_gradient;
