library verilog;
use verilog.vl_types.all;
entity tb_pts_sr_sv_unit is
end tb_pts_sr_sv_unit;
