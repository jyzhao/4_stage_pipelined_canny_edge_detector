library verilog;
use verilog.vl_types.all;
entity protein5_s is
    port(
        dbus0           : in     vl_logic_vector(4 downto 0);
        dout9           : in     vl_logic
    );
end protein5_s;
