library verilog;
use verilog.vl_types.all;
entity tb_sensor_s is
end tb_sensor_s;
